`timescale 1 ns / 100 ps
module lfsr128 
    (
    clk,
    resetn,
    clear,
    enable,
    load,
    din,
    q
    );
    
input               clk;
input               resetn;
input               clear;
input               enable;
input               load;
input   [127:0]     din;
output  [127:0]     q;  

reg     [127:0]     q;

always @ (posedge clk or negedge resetn) begin
    if (resetn==0) begin
        q[127:0] <= 128'h0123456789abcdeffedcba9876543210;
    end
    else begin
        if (clear == 1)         
            q[127:0] <= 128'h0123456789abcdeffedcba9876543210;
        else if (load == 1)
            q[127:0] <= din;
        else if (enable == 1)
        begin
            q[0] <= q[97] ^ q[100] ^ 1 ;
            q[1] <= q[98] ^ q[101] ^ 1 ;
            q[2] <= q[99] ^ q[102] ^ 1 ;
            q[3] <= q[100] ^ q[103] ^ 1 ;
            q[4] <= q[101] ^ q[104] ^ 1 ;
            q[5] <= q[102] ^ q[105] ^ 1 ;
            q[6] <= q[103] ^ q[106] ^ 1 ;
            q[7] <= q[104] ^ q[107] ^ 1 ;
            q[8] <= q[105] ^ q[108] ^ 1 ;
            q[9] <= q[106] ^ q[109] ^ 1 ;
            q[10] <= q[107] ^ q[110] ^ 1 ;
            q[11] <= q[108] ^ q[111] ^ 1 ;
            q[12] <= q[109] ^ q[112] ^ 1 ;
            q[13] <= q[110] ^ q[113] ^ 1 ;
            q[14] <= q[111] ^ q[114] ^ 1 ;
            q[15] <= q[112] ^ q[115] ^ 1 ;
            q[16] <= q[113] ^ q[116] ^ 1 ;
            q[17] <= q[114] ^ q[117] ^ 1 ;
            q[18] <= q[115] ^ q[118] ^ 1 ;
            q[19] <= q[116] ^ q[119] ^ 1 ;
            q[20] <= q[117] ^ q[120] ^ 1 ;
            q[21] <= q[118] ^ q[121] ^ 1 ;
            q[22] <= q[119] ^ q[122] ^ 1 ;
            q[23] <= q[120] ^ q[123] ^ 1 ;
            q[24] <= q[121] ^ q[124] ^ 1 ;
            q[25] <= q[122] ^ q[125] ^ 1 ;
            q[26] <= q[123] ^ q[126] ^ 1 ;
            q[27] <= q[124] ^ q[127] ^ 1 ;
            q[28] <= q[97] ^ q[100] ^ q[125] ^ 1 ;
            q[29] <= q[98] ^ q[101] ^ q[126] ^ 1 ;
            q[30] <= q[99] ^ q[102] ^ q[127] ^ 1 ;
            q[31] <= q[97] ^ q[103] ^ 1 ;
            q[32] <= q[98] ^ q[104] ^ 1 ;
            q[33] <= q[99] ^ q[105] ^ 1 ;
            q[34] <= q[100] ^ q[106] ^ 1 ;
            q[35] <= q[101] ^ q[107] ^ 1 ;
            q[36] <= q[102] ^ q[108] ^ 1 ;
            q[37] <= q[103] ^ q[109] ^ 1 ;
            q[38] <= q[104] ^ q[110] ^ 1 ;
            q[39] <= q[105] ^ q[111] ^ 1 ;
            q[40] <= q[106] ^ q[112] ^ 1 ;
            q[41] <= q[107] ^ q[113] ^ 1 ;
            q[42] <= q[108] ^ q[114] ^ 1 ;
            q[43] <= q[109] ^ q[115] ^ 1 ;
            q[44] <= q[110] ^ q[116] ^ 1 ;
            q[45] <= q[111] ^ q[117] ^ 1 ;
            q[46] <= q[112] ^ q[118] ^ 1 ;
            q[47] <= q[113] ^ q[119] ^ 1 ;
            q[48] <= q[114] ^ q[120] ^ 1 ;
            q[49] <= q[115] ^ q[121] ^ 1 ;
            q[50] <= q[116] ^ q[122] ^ 1 ;
            q[51] <= q[117] ^ q[123] ^ 1 ;
            q[52] <= q[118] ^ q[124] ^ 1 ;
            q[53] <= q[119] ^ q[125] ^ 1 ;
            q[54] <= q[120] ^ q[126] ^ 1 ;
            q[55] <= q[121] ^ q[127] ^ 1 ;
            q[56] <= q[97] ^ q[100] ^ q[122] ^ 1 ;
            q[57] <= q[98] ^ q[101] ^ q[123] ^ 1 ;
            q[58] <= q[99] ^ q[102] ^ q[124] ^ 1 ;
            q[59] <= q[100] ^ q[103] ^ q[125] ^ 1 ;
            q[60] <= q[101] ^ q[104] ^ q[126] ^ 1 ;
            q[61] <= q[102] ^ q[105] ^ q[127] ^ 1 ;
            q[62] <= q[97] ^ q[100] ^ q[103] ^ q[106] ^ 1 ;
            q[63] <= q[98] ^ q[101] ^ q[104] ^ q[107] ^ 1 ;
            q[64] <= q[99] ^ q[102] ^ q[105] ^ q[108] ^ 1 ;
            q[65] <= q[100] ^ q[103] ^ q[106] ^ q[109] ^ 1 ;
            q[66] <= q[101] ^ q[104] ^ q[107] ^ q[110] ^ 1 ;
            q[67] <= q[102] ^ q[105] ^ q[108] ^ q[111] ^ 1 ;
            q[68] <= q[103] ^ q[106] ^ q[109] ^ q[112] ^ 1 ;
            q[69] <= q[104] ^ q[107] ^ q[110] ^ q[113] ^ 1 ;
            q[70] <= q[105] ^ q[108] ^ q[111] ^ q[114] ^ 1 ;
            q[71] <= q[106] ^ q[109] ^ q[112] ^ q[115] ^ 1 ;
            q[72] <= q[107] ^ q[110] ^ q[113] ^ q[116] ^ 1 ;
            q[73] <= q[108] ^ q[111] ^ q[114] ^ q[117] ^ 1 ;
            q[74] <= q[109] ^ q[112] ^ q[115] ^ q[118] ^ 1 ;
            q[75] <= q[110] ^ q[113] ^ q[116] ^ q[119] ^ 1 ;
            q[76] <= q[111] ^ q[114] ^ q[117] ^ q[120] ^ 1 ;
            q[77] <= q[112] ^ q[115] ^ q[118] ^ q[121] ^ 1 ;
            q[78] <= q[113] ^ q[116] ^ q[119] ^ q[122] ^ 1 ;
            q[79] <= q[114] ^ q[117] ^ q[120] ^ q[123] ^ 1 ;
            q[80] <= q[115] ^ q[118] ^ q[121] ^ q[124] ^ 1 ;
            q[81] <= q[116] ^ q[119] ^ q[122] ^ q[125] ^ 1 ;
            q[82] <= q[117] ^ q[120] ^ q[123] ^ q[126] ^ 1 ;
            q[83] <= q[118] ^ q[121] ^ q[124] ^ q[127] ^ 1 ;
            q[84] <= q[97] ^ q[100] ^ q[119] ^ q[122] ^ q[125] ^ 1 ;
            q[85] <= q[98] ^ q[101] ^ q[120] ^ q[123] ^ q[126] ^ 1 ;
            q[86] <= q[99] ^ q[102] ^ q[121] ^ q[124] ^ q[127] ^ 1 ;
            q[87] <= q[97] ^ q[103] ^ q[122] ^ q[125] ^ 1 ;
            q[88] <= q[98] ^ q[104] ^ q[123] ^ q[126] ^ 1 ;
            q[89] <= q[99] ^ q[105] ^ q[124] ^ q[127] ^ 1 ;
            q[90] <= q[97] ^ q[106] ^ q[125] ^ 1 ;
            q[91] <= q[98] ^ q[107] ^ q[126] ^ 1 ;
            q[92] <= q[99] ^ q[108] ^ q[127] ^ 1 ;
            q[93] <= q[97] ^ q[109] ^ 1 ;
            q[94] <= q[98] ^ q[110] ^ 1 ;
            q[95] <= q[99] ^ q[111] ^ 1 ;
            q[96] <= q[100] ^ q[112] ^ 1 ;
            q[97] <= q[101] ^ q[113] ^ 1 ;
            q[98] <= q[102] ^ q[114] ^ 1 ;
            q[99] <= q[103] ^ q[115] ^ 1 ;
            q[100] <= q[104] ^ q[116] ^ 1 ;
            q[101] <= q[105] ^ q[117] ^ 1 ;
            q[102] <= q[106] ^ q[118] ^ 1 ;
            q[103] <= q[107] ^ q[119] ^ 1 ;
            q[104] <= q[108] ^ q[120] ^ 1 ;
            q[105] <= q[109] ^ q[121] ^ 1 ;
            q[106] <= q[110] ^ q[122] ^ 1 ;
            q[107] <= q[111] ^ q[123] ^ 1 ;
            q[108] <= q[112] ^ q[124] ^ 1 ;
            q[109] <= q[113] ^ q[125] ^ 1 ;
            q[110] <= q[114] ^ q[126] ^ 1 ;
            q[111] <= q[115] ^ q[127] ^ 1 ;
            q[112] <= q[97] ^ q[100] ^ q[116] ^ 1 ;
            q[113] <= q[98] ^ q[101] ^ q[117] ^ 1 ;
            q[114] <= q[99] ^ q[102] ^ q[118] ^ 1 ;
            q[115] <= q[100] ^ q[103] ^ q[119] ^ 1 ;
            q[116] <= q[101] ^ q[104] ^ q[120] ^ 1 ;
            q[117] <= q[102] ^ q[105] ^ q[121] ^ 1 ;
            q[118] <= q[103] ^ q[106] ^ q[122] ^ 1 ;
            q[119] <= q[104] ^ q[107] ^ q[123] ^ 1 ;
            q[120] <= q[105] ^ q[108] ^ q[124] ^ 1 ;
            q[121] <= q[106] ^ q[109] ^ q[125] ^ 1 ;
            q[122] <= q[107] ^ q[110] ^ q[126] ^ 1 ;
            q[123] <= q[108] ^ q[111] ^ q[127] ^ 1 ;
            q[124] <= q[97] ^ q[100] ^ q[109] ^ q[112] ^ 1 ;
            q[125] <= q[98] ^ q[101] ^ q[110] ^ q[113] ^ 1 ;
            q[126] <= q[99] ^ q[102] ^ q[111] ^ q[114] ^ 1 ;
            q[127] <= q[100] ^ q[103] ^ q[112] ^ q[115] ^ 1 ;
        end
    end
end

endmodule
